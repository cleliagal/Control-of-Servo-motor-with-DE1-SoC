library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- 
--entity clk64kHz is
--    Port (
--        clk    : in  STD_LOGIC;
--        reset  : in  STD_LOGIC;
--        clk_out: out STD_LOGIC
--    );
--end clk64kHz;
-- 
--architecture Behavioral of clk64kHz is
--    signal temporal: STD_LOGIC;
--    signal counter : integer range 0 to 780 := 0;
--begin
--    freq_divider: process (reset, clk) begin
--        if (reset = '1') then
--            temporal <= '0';
--            counter  <= 0;
--        elsif rising_edge(clk) then
--            if (counter = 780) then
--                temporal <= NOT(temporal);
--                counter  <= 0;
--            else
--                counter <= counter + 1;
--            end if;
--        end if;
--    end process;
-- 
--    clk_out <= temporal;
--end Behavioral;

--
--
--
--entity servo_pwm is
--    PORT (
--        clk   : IN  STD_LOGIC;
--        reset : IN  STD_LOGIC;
--        pos   : IN  STD_LOGIC_VECTOR(6 downto 0);
--        servo : OUT STD_LOGIC
--    );
--end servo_pwm;
--
--architecture Behavioral of servo_pwm is
--    -- Counter, from 0 to 1279.
--    signal cnt : unsigned(10 downto 0);
--    -- Temporal signal used to generate the PWM pulse.
--    signal pwmi: unsigned(7 downto 0);
--begin
--    -- Minimum value should be 0.5ms.
--    pwmi <= unsigned('0' & pos) + 32;
--    -- Counter process, from 0 to 1279.
--    counter: process (reset, clk) begin
--        if (reset = '1') then
--            cnt <= (others => '0');
--        elsif rising_edge(clk) then
--            if (cnt = 1279) then
--                cnt <= (others => '0');
--            else
--                cnt <= cnt + 1;
--            end if;
--        end if;
--    end process;
--    -- Output signal for the servomotor.
--    servo <= '1' when (cnt < pwmi) else '0';
--end Behavioral;
--
--

--
--
--
--entity servo_pwm_clk64kHz is
--    PORT(
--        clk  : IN  STD_LOGIC;
--        reset: IN  STD_LOGIC;
--        pos  : IN  STD_LOGIC_VECTOR(6 downto 0);
--        servo: OUT STD_LOGIC
--    );
--end servo_pwm_clk64kHz;
--
--architecture Behavioral of servo_pwm_clk64kHz is
--    COMPONENT clk64kHz
--        PORT(
--            clk    : in  STD_LOGIC;
--            reset  : in  STD_LOGIC;
--            clk_out: out STD_LOGIC
--        );
--    END COMPONENT;
--    
--    COMPONENT servo_pwm
--        PORT (
--            clk   : IN  STD_LOGIC;
--            reset : IN  STD_LOGIC;
--            pos   : IN  STD_LOGIC_VECTOR(6 downto 0);
--            servo : OUT STD_LOGIC
--        );
--    END COMPONENT;
--    
--    signal clk_out : STD_LOGIC := '0';
--	 
--	 
--begin
--    clk64kHz_map: clk64kHz PORT MAP(
--        clk => clk, 
--		  reset => reset, 
--		  clk_out => clk
--    );
--    
--    servo_pwm_map: servo_pwm PORT MAP(
--        clk_out => clk_out,
--		  reset => reset,
--		  pos => pos,
--		  servo => servo
--    );
--end Behavioral;
--
--
--
--
--
--
--ENTITY servo_pwm_clk64kHz_tb IS
--END servo_pwm_clk64kHz_tb;
-- 
--ARCHITECTURE behavior OF servo_pwm_clk64kHz_tb IS
--    -- Unit under test.
--    COMPONENT servo_pwm_clk64kHz
--        PORT(
--            clk   : IN  std_logic;
--            reset : IN  std_logic;
--            pos   : IN  std_logic_vector(6 downto 0);
--            servo : OUT std_logic
--        );
--    END COMPONENT;
--
--    -- Inputs.
--    signal clk  : std_logic := '0';
--    signal reset: std_logic := '0';
--    signal pos  : std_logic_vector(6 downto 0) := (others => '0');
--    -- Outputs.
--    signal servo : std_logic;
--    -- Clock definition.
--    constant clk_period : time := 10 ns;
--BEGIN
--    -- Instance of the unit under test.
--    uut: servo_pwm_clk64kHz PORT MAP (
--        clk => clk,
--        reset => reset,
--        pos => pos,
--        servo => servo
--    );
--
--   -- Definition of the clock process.
--   clk_process :process begin
--        clk <= '0';
--        wait for clk_period/2;
--        clk <= '1';
--        wait for clk_period/2;
--   end process;
-- 
--    -- Stimuli process.
--    stimuli: process begin
--        reset <= '1';
--        wait for 50 ns;
--        reset <= '0';
--        wait for 50 ns;
--        pos <= "0000000";
--        wait for 20 ms;
--        pos <= "0101000";
--        wait for 20 ms;
--        pos <= "1010000";
--        wait for 20 ms;
--        pos <= "1111000";
--        wait for 20 ms;
--        pos <= "1111111";
--        wait;
--    end process;
--END;